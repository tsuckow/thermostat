package lcd;

   typedef struct
   {
      logic [7:0] r;
      logic [7:0] g;
      logic [7:0] b;
   } color;

endpackage

